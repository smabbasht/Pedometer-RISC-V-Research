module pedometer(

);
    
    
endmodule