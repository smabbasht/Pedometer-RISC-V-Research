`include "node.v";

module ExBlock();
    input  [9:0] A, B;  // Our inputs X and Y
    input  [2:0] funct; // Determines the type of instructions
    output step;        // Our Final Boolean Output

endmodule